XlxV64EB    17ed     730�HGU���Et+�u�{�v�|M
o���3�����/��n��غ&��M �\��C�q!�5� �o���g��}��1R$�'�0K�E6�V3(o�S8 ~'63�>Z`�z��(��̑�`Nwu�a�y�b@X:������ O*56Y����.���GF��D�W�tA��o�)��=�[I;m��J��E����{�OήЬ�T��F���
>}�X���S���M�t?������X�6���AI4��
ln��at�q�.�f�Ҫ�(���|��äO��f��
*;v��=������|��������5�q�]������e5c.�?��I�hfJ?_Z��Sg(}�H�U��:t�+nߠ4~^M@���ť]���;��!AvQ9ԥ�EͲ���������GL�&#ˎ$Zq	'�ެ��ѠڜV�l�^�
�5�E�
�ԩ@��8��K�#=�͉�t��i�����yl��_��6�;&�����QHJ�a�����%�sC���W==x�������ÓM�'#\С���?�M���V�'��O{V��=HX�����8�W��3c"��9g<�/?�v�	\��U��x�}
P�������$u΍zq\ �o��J���d��L)Q }p�7�;�'��N�>�h򉎣ԲJ��?'7ψC�����֣?f 5�Zb��s" J���(�f0Z���/�>��Hˀ��'&�����齝����	fa���<E&w�|�vm��c[��~����H˟Iq�n������0��%�K�!�d�0�뗽����}��������5=/�V�ۺ	v�U�|��+���vX҆��<k�O��k���	b�n����c��m�����Jh^�}���H��xWG��a~�7���Nb�~*h��QÌ�-�zݨJ*|�&�o��@�_���z-��d>C�;��}Nm]	Ƌ����Hl�C �����TH��R����W&�v {iPB�ot����d�m����g��8�L�=�oz��ú�;o�~��mv ��Y)���8�\NÚ[�Z��2_����H���L(#Ƞ�])���] !�kq��m2��q,~�MH�[��t}$�"�?��H_i��a��1������PWOy/S��cp�z�"���@�#Sn��dVȟsMŖ�$%��L�x�$Gy*�3]0l��F���0��`#/���:p;�j;φ;[���v�-~���X�y9z�}9E^�|U��Q��Ϩ�7\{eԙ�
���s�/�HQ��=;&3F���q�o��&zw�E�w����b��Vj �u��H\c��i�ڦod����G��Q��n�zȫJڭ�J�!��ǮIW�H��%��.��]h|�L󴅢��� 8��/c��}���ϗ�u$�c���b?�I��5/	�Ww(d6#�AsA��
��8��4�C}�V�7�=Z]67�G��M0D'b6��S���i�,f�+Ȥ�ca �R��}�@�iy�[�ᓦJb�\�@��tmyn��u@o�U�^�Pi����xE�W�Dq'��K@�c�_3�P|	��퓵�ئ��H�X& 0L�qxe�,!��DhR�i,7�'E�@�n�=r>h�k>A�S,����:쐞�Ҙ��Q�ر�
P���&�#�n����}m��?&7id��K򏭶�|6<�JU�����̑1r�0��r������zL��`���6���n;���P�dZ!�B�k��"u���;Λ\�9ըe��N����"ɯ��S�i�����Uj�qxh�Z8�͋�6�~���J�8@/�T����gi��m�M��@�