XlxV64EB     e36     6d0������1qa��K�V\Į���4gی�z,�i��9ĠnM���}���K��*B�@���p��_��V�)y���-�O;��+���]���6m!������m�}��!c����������'�sO�������ӳ�'�	#ViP�2L�6j��v���)m�Σ��;GнI"OYK��;J
ᴐ-�	�IP��PL;H����w��z*V����.][�y�)��ח4r¸�K�^�yc�ͳ,KԹ���܃IpŘ6��$����	-��t�x�0��͕n�hv����m_��'�ʺ�]�#k�ӿ<,@z�mY��G:/���v�h�z�%��AI�3]wI<����*`S���y�E��Ь����F�I�x�XM��鏇�I�'>���T����zvɢ��biR��~`�,�=��u�ZR����4�H�h�׷)c���c�'0��Vw�-&�s-�i�-����&TsK'/����@�s_�,s��Ւ2��z3*Qa�K�kBE�	$L� )sˮ��a��:�*Em0�Ä���]�{J���T0��U��,,��,G��;uM��w��������(�=���ڦ`Վ�hWO�\���迥:j��f?P�U	�~6�G��������G��-T��'��,_�``�#9ȡ.�.q����FJ�L ��[1T^���W��í����N�V����;� ��)��N�V�PE�ord�����������h{���ӟ���1��C��7`ܟ�Y\;5eD�{�M+A�9q����EJH�Ocq�x��PT����(�4�l���f[M��w�r�IN�f6����A-D��Ңf����V姡�Y[����Ŵ��WÎ5֦ϟ��ܫj6CҦ��w��is6����	�k�W��U{x����,�vl���/��C�1f=˺+HH|v�GY�[��hiTm��i�5dJ�T������[��vL áo�i�W�M �ʏG+��~nl�!�Uz&���e��T����+�_$b&G
�ښkw�+��t����M��޹m������`��8!��?LY2Z���:DXTgt�����o����i��������t�t��МA��o&ĈJȀbCI�ϥ6|w|����顡��>O�zpn�� "������	���4R�܀��[I�t(G4goV.�xqAny��~��z}��OD�ja��dp�V:k0{�x���Y}�>�ũ��d��<ٖ`e���, ��T�]����"/�:N|szy:(9�M��[q�N�e����c�Cc�(BᶯcR�˘��!�.z��� ���[#÷ejtP��ic쐉j�4I1/kS�tt����lٴew�f������jr�e�H�a�G}��l1굽��l�%>�`��3��
��������5q�`l�&��y��^�7:�؉
У3t�)�)���^�g�tv�Iyb��� )[w��24����Is�B���Y#6e��DL�Q�E��X�O��+��T����	�O�����r�#&����uf��ĸ���!ƬXQ���}�eUu]�����-�"���:�H�Ep��3[�q��_�6�%jV�����c����M/�%A�
yܿ���l��Q	k��Zo0�٦-�?�!]S�!�8[\>ϊ~�j�k���U���E�G�+2Zt�h��^�A���IL��R�L�ƃ|E[���y���b�?V@+�ea}��+ʳ���j%:���z�