XlxV64EB    fa00    30f0�%���B����#�/���	����n�d�1y|r ��|�VK�
fr�j�@8=��̏?%{S�(����8���`�����0�2���>��kӍ �NdE=�*��'	��������l� F;K�����T�L�V����&�j�0��ePPxC�<�=�p�se�r5��M�)��Lw=��w��h®�CBf�U��g��Q�N��rߝM�;�����hi�X�X��e�K�v������h�l��,;�ܔ�y��@u�$qu�����Ob�2$0�vsV�v���}Ͷ�xb I�\F��ޣ]��,��V�����w�Y��$����<=�z����g�����q�U��A�ޝ�{���Z�����N�@Mh ܥ��u�a�S�X�RT
��:�}�h3@��%HTN@�[�.���َ��e/%�+��>/7�"Y���e*�(z�ʘ��1��<Ö�'�7���B�e�2L2T|�K��-���nߺa��ЋL���/����Ց8��r"!����K9���K��'t^�����0�Y��F����B���x����̽����_�zN��K4�#�WG��Lg�k)���>�0O��1�=�:Ƅ��XV�l燎M~��v���W[[�b*l>ştRZ'"�!N��@��p`	�?��\�Z.��G-t����?�W����ӧ�^E>��@&�����2�k k�F[m6���֐�}6�Z�
��<xF��q�/�Xj�CV�f��K�g��4�/O:���)��Z�Ĝi�@����`no�Q﹄(ݟ��k��{B�@)a��TW�1g����	\�Y�І&�h4�[��c�|l?���E���|��&�ow(w�οk��؊��`0�b�ǋ���(��Z)�<�]�< �W�ӑ��,&b�.�.#����_ۥ�/* 2x�4�|Β1ܦ�����M���J�1�H�O����eg�b�4u�!Th�;9����y�'Q��94���y@�I�Q˟.�0'��?��-��% x�S��LSo�G?�`�}RBF	{��C��M�VI���7<yD�[u�|�Z��F�$��
�"�:�r௭h��i��ω��p+�#;qXu��'�Y_A�G�+O�M��o�?��{���n����ѻ��Z�yp�9ā�:�Lz�9�5�u{�Z��p�1�yN�vK[s%e��!�A�W����o�t�օ	�$�J�ܼ�>�.��N�5���N�̱�/��<<*�t�o����ō��JOx����)��z��>���9D>��r���VжD�Ki�$� �=�r�C#6RE͉�:�3�)i���O׻��_�ͨH�O�5?eٙ��imB��h������7�s��x�aO�h�}��bZؼA�md0F��'Cb6c�ٷa�qx��iy�:�Q@��Q=̲�`�$�יc��:���Yo��b��I� ��,8)��xi�X3ۂ�S[�u�����8�3\)����v��O�
#';4ǰ�[K�i���
��a0�}}��|2J?�Wɪ,/����L����M%��㸜����s�?��;f�7�o뙆���Q{w����C;��N��*�,�1�@���0l���k	���f3e:L�tB#^��%�ۊ�sV�PU`@	}IJ]r�|2�B�e��ݑӐnH�K��
]�ݍV����Lf���q�7��	�xB�<9��a�sGg����fX��f�WVJXDP�4�B��8YH�t?w�_�0�͌��[���a�7��RASފ��ğN���e�P���^yce%�)��6�����A�,P~�X�܁ĳ�\����k����YMG	|��S
 GbyE��/.�{�p���h,A��-��~N�
���"?������[z�b1S�NTd�ֻ�����;�E��w,���P���riB �N��C�b�e)i�7�_�-�>����B���7�Ibb��^1���Y�8�/r����`�b|cAb�g�q��v���j�[)�P� +�ԝ�j�$��m��}�`0/�X!��Wa@J?����&�X$@�qA��6�/����+I�bo�K�`<��)���H�����������ς�r��NهS	=5̦ظOB)d����^������Tc��|V��n�6��H�Q���|����}>#ri9��`��k^<z7_;2�ɖ�@��l�O!b�:��5�EF���
�ʓ��W���bL�?@�FJ}ܳciK��l!''�<��'��W6{�u%�G��LbZ�Wx��N�� �voO!n�3�𼏡�U� �K%� ��~��F*�Ȱ� ɒ�O>Nh㜨4-��:D-�K:���Νw`�h/��K�6o;bK/�ÑI�.�A�Y�҉w�����t�(҃�LK��x���:K��=B4XE����f����w����0�p��,'\|�1���UO���8
^5y#$��gY�K���^[ZDyϫ�#K����~�e�f�e��i(˵i��٣�q�e�s�k87:�;�V��,�M�rz�Rs5AG*F������i4�FsT�N2�	U3�]�=��<j��/@�s�p,y�b��`�#���A�J�n
vc�ُ��_b&�ac>��-[��� (�2Q��|sŖԇ��(��X�*�V7=?N�0K�ܧ-���r��;��j�� m��`O5�D:X�U��O�M�T��A�Y{�i�����o�K+7��E�ܐ����f��ܑj��1��y����K�]�^_V���x�3�X�I��z�~�Ә�	�L��${!n����*mx�Z֎(:�T��H��	���i����@��h'��#X����0�H)f5��]������Սi�ir4����/�-�h%��������smVƭ�|��2Y팍��*��~��f���-	�b70t�,��L�"!Ge��e�>��%>��U���)�ؓ��r��	�[2Sw5}�jZn�E�9kH���h�'�C3��<w��1&D=DfE�$ �M��s�uf=C}^ζx��%  U������8E��#}���`�{� �|��k"��kf��)_*?����t��/�ܣn�ȯ8�ԣ�C*Rh�����CY8\:��'n|�U[\��{��_�:fy������ƜF��rzjD��-*7��է&��=E�$S�L���V�k2r��tn���'?-o��ђV-�2�	iQ�t0<�pD�Q�;���=�+���˨��W�uhL���=��U��:^�~�Sru-#�e���m��ݕ��i�⊇�xS�QM"�Xjq&�;ڊi�9�^`�r�m�����lk��S�WS8Tr�D�@����3�o۷&yf�_�d�#��M�Ch�4�%v�Jԉ�����V+Z��/� �g�ɾ���2�.�hY��D���qj��39t~�4g=/q�b��&/���QOK�%j���&�t��:�J�<E*椤j?E�T8v&��h{u�?�T3n��!n�&>i~��H;�0H�x����oi"�Y׼�.B_���>���!}4{��e0�o<��/��Q����k �0-�d�Ddb�|0�Q�q���A�*�Opק	���o��	#�A��gy��[8�����e_[]A��ߛ���s�q.^i
kq@���|_�LJ};��sv�wLB�{�*JF�(�|�$%o��T���'b4�I6�+�Ԟ'��Jk�CA�����l�K�OΙ^B�x���ȅ%M��Kv���ζ�K7�m��`A���ǔ����.P}��Vp��uN&�)��_D������>;�$ޠy�q��d���د�+���%��3��2@��0�Ez��ř��Ɯ5'��p�������R쥊�'��=��0��u���w�^{���A�����dG�\�b�J�?J�9�d���*l�ևt�m���^��_�%\�_��+�֬;�K���\)6�
��v����;��F��ۑ���G�,��%A�K�?��[�M�3s�*%�p�+�SЮ�y����݆3�*���ˏ]G�7�7{&`�Hl�~�޿Q��G%	$����@����U.(�v8�ҚA�2��r$�x��Y�µb6��
.�!�	�� �՞�t�i0W*�J���N��������М�zwb"����4����k�KVe��1��!-��u̲?��*8�%W�o�&t{�枷Ȩ�k+�x`RRJoD�Q��^�L-��
���q�">	�!�_�?�Q��<��7�yuR�֮�)���X�4�:���4���%���ٳ��6�xGJ�o�GP�j�������P m8���j��Aq+R�H&�l�OoOSt����jQ��r������>Rk�Ɩ�➾����T�V'
Yz2r\��o�7�wu����֦��{F������v�̤�0����C�{	���t���$�D*=~ic%b2j:..۱����m��r�.ˢ!��d]��y8).L��_VH�0���;cm�����W�����{ #�{��_�o�_�o+�#�s*�t��u���PT.�P�����(j�'��+�}��gp�)8R���$�I�%�D�?�P�Y-���9?*����$^��k�%�SL+Rɲj=&�{k�o]�C8����x�j��pw��Ϧ��³ݳF��4��5.���w�C\ݟ��Uv��>�O[�
(,u��yj�R�x�E�6��9����=���j6���D� [	���s5k#RJ��x��s��He
�_�+�^k�U�Ё��ٛO�TƤ���8�و� �yۤ�fv���&�q���`��M�$��}������76ǰ���Fu�H���i80��Q2�4��[�atC��D!A	6���#@�I��bc�F���U���]ғ�4��5F.����ў��%�Q�F���.����GgH Π<���	u
��{�G��uH�T0ږǶB��6�H�a����K4��<��<��z1�ȁR2�*o�u���K�[���I\�h�h�l�b$�r[U�=�1H|�}jMWd`�4�Rk�Aj�\�.<�=���m���?Z~j�%�Ǟ?��z�b�e!��Ti�VRk[�P,4؈c�uvHdGnr��0�n�_��Ckc8�h��_L��g���\�Pv3@����%�d���&����Ih���J��$Z��S����"j�4�H�	� ��Iz�JO�����n�l�"3�>��uԏ�z���V�w�$�	C���L_W�Ԣ�W���N��x��#e�l��O�쩭oP�Q{���������_��M+4�j�=�/�/���`�S�cgak��������D���N�����E��AA{Ĥ�Ys�^��=�?��L���CM;����0F���j�d���ho�e���p
J������u�n��Dv(��9����B����U��:��wG���r��JR�^|��E�Da���QmI:Vb���\�,\�	����W_�X	?!�Q�
�K���q��*�68g\S����y�<��J}����s7�|@R2�1R!b�Q�b�$���=9̈́t��v���^�N�jq�
_$ɨ���n��9v�(�]��q{�@v#�;H�Y�*�+�#fՎ!|f�	#����w���~Լ�G�u�u1�FuM�}Dl��������z�
.Lg5Qxg�����=#.�Xi(��}��5�� ae<����j>��f�V���</��=�l�8}@�)�J^lZ����[f�g�6piq{S���`Z$O��%���c}�x���^i�7tԀ��'�b������2�ON�M�-{Q�_��o�h���e[�%x��_o,�̩���sB��t��* a�?�'���Q�7��s�,kKԚ�J�.$\�d��t���U82�F�&�z�]d�Hg���`�0J�H��^Rd/��R4^����ό����¿�+Ү�q�p���Au(4�(K�A�+h�H_�q7upOD���pv.\ hl�v��95�ݧ�L�T~���%�
T��(rq=�ƈ�]6������i�K4��WJ�_��� ]�@���ls��m��4�j�d��G6@/	�>�aZojH{��X~ߥ�!�����'����Gw�B˂��F�>��j֥��f6��kb!������i}%��o��k*�)@�+Le�+i�<�e�Y��E��-����<���ӻ���Q�-SZ���N��$q~�"��p��?R�Շ��L�z(� ̆��A^*x��X#�v�JF�"��V�V���L>�����/�.�|F)�H�4�=jU��VS��)~}��qs)�MP�z�#���ǢueZ��U��F�)��M��=g��E�d�P���g)rпq�	Z�\���w�u 6P	�L�5���!�7G��Ԩ�w�<д�vP�b �:�dԎ-��c��
&�7ͩ�5�����Q�*���|���$E�C�n;N��5�Y
�0Z��I����^
,�ls��,��;ߣ�:��c�p9W��N��B�`� i|�D&v�Q��p~v{�N5m��5}�@�y��9$:i����¥Q*{,����RݗH���qzn�?ƸH����^&7H.Yz&h�y�C��q^
�b���5��R�q�x�����i؀���.���[k�8���׃({��/�QE�i�#�v
r�`��`�魾4I8�R���̐2c��x!k�nY���+9,��V��ת��6"1����!��v�n���O�F�% O����i��9w�}Nq����G��<��I�)�Y��P�ʎd%�d?Ù"� ���d������A|>�ϖ�$��V>�:|�������@a�LC	O��+߀aH:,����^���ڈ��U��X��͖�J��"wd��%���&m-0R��֩�Shi 1Q�UԨ�$�F�r��^�|�#��Ʃ)�g�7�Ϯ��e�D�BS��܆��7(BH~�. ����u�Ule.�Dઁ�"��3�)ݥ����vBUA����l)� C��[��gQY����~��J�ٻ�Dw��0�	�X�>�P0�M���KF��p3��	��k���Y�gvZ��S�Q�"D���ןl@6�Z�k��ڪ�����pe-��`żF���s�p ��~�i�x�x9wL��.����ơ�\9���{Z����i�����M���i{Є���]x��p�Կ8�LP�^�Tt�џ�����h 5.����\�A�1��R������M�`�=�%���Ȣ�a}�*r\c�11����=��E��ΰ���Gx��>S��.��B�Ѥ�I��<�k��q�����BO�
|s.t;]7ި��&Xj94H���+&�(��2L�,�ͦ_�W�Ɉ���My�_��F�]Kw�ں�G�N^7ڠ:�JfB�Dʘ�=��o7�4k[�ϕ�`��"���ڳ�KY��kbd�w�H��vX](�U1�$Im�~�����jM:x`���D���$�­wL�x�qq����T�����!c�Ͼ��EK �E7"�����L��.m�0Wv�>�6K�>�6Q`��ųgƇV��Ӳ�O�!d�	����PnuQ粦nq��E�=��WC��4�Ԓ����w5{o���q���D�%����s#s����ɬuWG��h�Ӡ�#8���<�|`�T�����D^+I�p��lԭp�]��/77VTР;>������R�<w��K�^#����nH(�z���ɼ9�1������LA������܎ܥhs�N��l��M��y��W�}�Wބ�	���J&��ރ��t�������Y{/�ǉ&ݵ�A�s���>���7��d���C�kdU�%����L�͞%���_�r�[�'��>���~���Q#N�Z��?���P(	�,;l'�bA;;mK!:A��a���o�"Q�]�`dR
�Ԯݾy����5{Q܂����g����R_��!��Q:��������N�V��Q�h���+���M]�੖��VO[d��v��4~�U �T%�W-e�]y.��Q[*~�V;�v@\F�m\,�Z�,8f����x��1|�"�)p�����[`�Z�%S�\>H��8�$��m-�����5�0g���>"�k<��=������A�H-�*0��Oc=�I��,%�i� � ���������wJz��'�@��u�=�4��;qX��}�x�����M�h����s�i��q��N�P�S�i����u�ǲ�_����������	#�\����Wv�ۿ�����;(�5�?5ki����)~Z�2�[E�_�B[H�5���?���F�����L�s5d�k�1a�mΗv�����C��o����o�v��B]�Uk�D�F�n�M~�:��oʰ	}�)�O�VWnN�a�@��=���p5���uU<:��!�/�����H����3�c+}��n�t殘v�K~��3�:�ߧ�"'P��vE�]�BWx|���?��8q* �r�aπ�eť4�I����	v���i�����	b�!�3�-TS�)?6�w�y�Hy97�Vm�&��joR�j����.�	.���H�<��rݓ^�(��~�*�_k��n��˩̫�}��>?#췡��~���W���%��U�hnQ�9�务0����VT����o��gd�s��
g����m�+�C���~���b\�e���,��?�5�N56��B��Z%O���ƃ q������P~�k:es/��k����&2�� �q7T�j�|�$~9�MY�׸G��7B�[WC�
�>�9Z�|�;�d����F0�71��;�7y�c�$�c��-
e�T��s٪x�x�F�	��w��F�Hq������%���?�B�"m�lt�h�fs���j��I��s9��A��'��	�_���ư5�鿹ܺ$�a��U��P���|k<c_���w��e+���g�H�<���0��t?u?�=5W��D���ؤ_9<�b�/�� ��2x������2Z��.�3�
xy��]>ݨ�l��A������N|�a)\~�-{�/z��	`L�!Ό��[S(*�<���X�s�����)�y��%�������׸t��`�)�ÛC�6S��>Y��*��$�}�FΖe����c�=X��J�Ě1����04�z�o�Uy�-��d��Y �u-���e��-��x���p\�b-�f��Ջ�Ɯ�	�E���"�M �l��o�3�ա��Dc=�*���#�����Q�Rs< ���$��]+�jn��u}��D�Hr���A͘�� �b��S����HQ��6����G�n7��3s�	���]�_#4��8D�;��x�5�/�v?��.}��'2����ƭgA��]�4�p��k�� @�Ң���{c����=��]]
�h\�1��ZZQ�V�n'�z��c�Sn4���������~\c;;O�fA*t�}�h�����L�\������d|��Ϻ�Z.c�hZV̈i��f����S��L��T�sfqVu���9AH��39I��c�K93H�X�BԺ�B}4KVd��"���N.C�2����b]�"%��rx+�̨�
"dC ?�&�uф�����ט�t��P�|-=�#y��s��&秊)?��n�ޞ0�@\=U�m�0���)�D��7����%�l��$A��)}�~ÊQ1x
�l��0ᐢֻ(f��g�"�Q��I
��O$�I�n*VT(���?��h��&��?�n��� u��Mɀ�0r�sG����&>1 P��;�X>X��)���7UC�ݶ�����Ll��QɄ̷≯:�p,U��D/(�h
e*JԽT�����y$!�wN�r�?�Ԍ|
��Ħ�	嘦HG`d6c���t�mw�9����;,׵���UD0�h��2�}G�z�L�W����#8����ؕ�)���6R[�S���@��j�XvL�'d�ƎS
�}�<�N�E��m�K�%ݱ5\�b�ɳ�>��P�%V-�{�|�tyaY�μ�en�=���V!����*���r)/�Zp���pi�F:���j4<�w�*�S�j4��vUg��X3��eΏnS/_BF"�.j�fN��ѿ�H����b��6���������c��$���dzG��=b?/9�<�,�+p�������24��܏�[
Ҷ��r�^&�G\A�����e��e�qQ�M!����{k�f��0�7���n��՛qZ.\f�R����$��@�w#r%�1(�`6~]x��T�W�Ŝ���-y,�ۋ��MP���.//T�M�M�r89XHs������ !�3i.��0�a׻Dg��-��*4�;ޢ 	< RL(QT[l�J"���!�Ӳt��Ag)?-�Gq:��"o�P�r�8 ��2��\�uJP����ݣv:�_\ۭO_���}�7�C�ҢZ(� "����A nB;[�[ �M���`�VY��rNĿ�z�R�v����|?�&$�u�>4�hI:Lbc�-�"��l�C�~�d��n{��P�5�6�!�6R`��U����B(q�6�>p�k����Ad	B+�ł��M9�������)����RF	^�Mz����8�ۂ�~���Y._��x�P8��?�x�ڣ�$�4�u+V�e��P��ݕ@ �/^zG�|e,*oN��ʅGi.|Qc�A��ߖ�c�z�&jCP+�34�F�T�x�I����n�Oօ9K�>����������O3㚦�?{�^̜/aB׽�<��=����r�>���wK�#u� {�L�K��C�^5�����s߷#���4f�<�J;n�m�iBur���,��v�?.�D�I�R�-�?'fV����UX7�c\ӥ�RaU3���3�th�����;ad�xψxd�sh�
?����V�`��M�!r���]�<���1�R���3������`�Ԇ�1&�w!��}9�#*�,���%�z&������{6�m����!$��'V �Uɰ�q�_�O�XΟ]�!�+'�37��C?�tP���A�R&Z0w�:��%�=}'�+��;!S���[詇΀�o���@����M�_�3��C_5����i�Ძ��Ev<�7u���W2�.?1�2
�������
H&T���2��:�|�����l����s�� ��Sg��0�DO ۏ��ozG��R��!���B�u�4lwٖ�V�j/k~!�rwߜ�J�L8��b{�F�G�a�m�jO�	 L�@�W�����G�G�~e��iH(&�3�W���/�7V���ˬ��i�H��}��}��y�����ey.q��[�hn�:бL��w�&10�0}��'��������l퟈��D�'[}(�I�WyBzp>4�;L�AH3�lLZ"�[t�ʕG��zd�>�k�������*�xIb��Z���!���zص��h?��;u ��퇧SN�1��J9�H�j�����b�Fk;���^_;��~����V�_�a��s�Qx�5���s��隣�Ի?#�5�̲��W\ ��TE�ρ�X��z����b�/�����*�i?Hv�L�A��V�v�#��Y���c�]��r�r��.G�3����!"�D�@Y�'��/��K��j@�L�J{��r����Z��Ew^ /
0�Yg����tW��2콯Π�_?Up��|��̃��R[[�Aӷ�e����HkkQ�<:7JBe_�%�jx�ҍF��Ь��i� E��C�	��jB�<��^� ���&VM�B.�a�+f�f��mԤ���3��F�g��?����vPe�GdE��a+����] �Z	2��X�\�ۺQ���q�<��,��IM���y�M���$��@BM A�O`k��R�SR��#��H
�w7�OS 2���)U�֘�d�*m*w�D� �`�Z��3~�����;�)�,�ڻ�N%hN"�LE���DUȚ���v*	�����d��hfz����e�p$_���,�����H��mm�1�J:�tN��{/ ��&��w��B,��e.��)�ULn�|��rk�iI�/��n�����[Y�߮�Y�p	ٙ�l���A;2RU4Wt�罨i�����A@�����NJ��,T(Zj�y7rUd,X�����"��΁�H�0i�96�'��E9�{�u���KMGvZ�⸶�R�l��I;'w��X��k�hqt�H-������WUa�v&�� �W��*���+7����r���Š�<�;t7����C���֮a��W{j����B<�g���du�Ğj���9�+�J���I�b�en[+í�[�&fA#��=�I�X�rj#��W����dr��LIͱ�U�՚?gS��������XlxV64EB    ab23    1af0c����7�
4_�Pf��;������R2�Ub��t�n����II����1�_�N�=kr�=G�We��d�Ae�-e�b�����ڒ/*�~3��<:䆣��Z�z�[9�<H�~���m:����@b��y%i϶Z��ר讜�CZuu�7I�������FW���![�&��Qf�?��Q-��:<K��b�l-$4�H�O�P�U��R�F����:^�l�>4x��};,p����6��@IȝCa�DZ]y�p��w���͛���BzQ7��(����<��I�n�����]�
(��b>C���ey&l�ۗ	z���&������ϕOѸX0����!���퍺@6l���M�-c����X��)W���l5�z�k�Oŀ�T�*��\8I����eK�-*F[��齝����`�X>PLC�I�a���vȴR7� H5�pNԕ$�9j�-���$��g/�]�����ҟF̦5�o�5ic�rH�8�hs_J�.���ʦ_�0C�3����|�5��r4�8��������s��_�^��i$!RwT㫊��0:K��RB�%��t�(���;�{��aC�'�򇂂]�P���\ye�L
�n�L&�" �Ռ�/S/�ݑ���Ŧ�1Y,~�(^*�a�`.��'�Vh��D�g6�jәӾ�O�2o��B\��_Yxȉ���T/�d� l�B���*���z{uo+J�7�cZ
�'y�V)r�i�_�ֳ��y{�NS[���b��J�?*��M�����G�f�I���>��5��Iz�������-�"���%���'p�E��҇�I���OD��3���N�@�,g��f�S�ߣ�{bt>����#�]7�3�v"3��۷�~�;9��;���p�y�jK�os��(���&����衍,��F��,���A{���ο��d����a��6�X��h����Y9��N�]ګ�c�����:�U(�'
�/��RI"��M������Z烴��Z����ʗs�u�ӢcWE�],��gV�e�.�boo�ڷ�6Y.-� z����h���P�O=�؈�� �UOmO��3)��
�7��=��<N��s�wl�JgI�z1��3�E��C�q�A;X�·�����\�y{~����I�m�!�$���j\y<<)G�Q�^P��i����&�,Y�$��x�m��7j�xh���k�ӎ"��Ј�>��Y����쒬�ѹ5�E�e�*f{�Lҽ�_ϱ�KZP��Í�ޝ�fN[1D9�h@Um
���$+�w<�
�b�z�;,>�=�λ"����<{�뺬^wܣ�[{��b��,��]��j�6r��uHଟ?l�ae�H��ja�W�V#��̧I�lW�b1�G�Y�R��'ֵ{k�D�'";-si �Zn�
����o#��{��:�N�<[�`~�y%���m0�^�6OR�&��d��/S��u������A0�w��iB��W��l���FD��I��%���W�♮WM���@�_E"�c?���h�aiUpFk�k ����I�(�=x��\�H ��\r����G���04�)%��\>��p~F�Ⱡ��s����S2,]����ʽ�mN��5x {`S�^M+�xrh�@*��f�K����DU��5 �]L��7<�K���J�sjWm�1*�`é���JF��0���l{���ӘA|B�󴧟��R�wIu�����X�OFj�m/�߿o�%%]�]_�o�aV��́�����sU&�9���c�V.7
~v�W�+#;\� 	����k>�}4?��:��wA���o3�!�sT[QJ1�[��lo;��Tܒ�L���Y���)7����!)��D'}JJ)�`��;�K� %P���D�\3�K>�{����)U�H`ٵ(3�ʤ��.n���X�~�9aEU`�����*b��BV��'W+�b+QH��.����0bkJ��|�Tۜq��X��\2�)d:��v��7�6A�L#�6�!���u������t��/���	KJ2��m~9)�\�*�Q�\p*#���)|���I���Ȧi�aURx;Il��<G^���ɽ��`�[m]�?���I/�tc��ůR'����*�rzC����Ȳw��K�jx.�����@Ò��|T@��q5����z����z�4?~f��<lm�#�+�J��[�[��L����Z�姘�C	a��/��Zc�p
g�M���ꩤ�;�d���2L+�	BcQ`;��a��7ċ\ɏ�6WZ�If�cr�2Y$���
<v�R�2O	���/����PC��	��~*)�d���R�$࿟E���W��b���	�f'r����v2�F��J���Fx>yX��i�4E�����5�`���%�}�����>/��~�j�?W}��©�l=Y;�İ�e��~(#�V�n�$���� !8� ��?��cxN�~]˿��>�x>����yU��i�R�>��UQe��Qd�{5�9�k��ގ���ڬ@t�Q���~�@/�DU���
["WҲ{l�#�y��I���A���o��ᑦA���%��B�2�X�8jR/���9�8���3Q��s�l w���P�}�K�^����Q�����0R󜘛f��H~X*�q;�A���=L�Z�R��ѝ+���	ISf�֏�k\��2�������ױ���̐���h��p"_l7j�T�3zfL<	?a�o�"��Q	��T�UGAK��Z�2�r��w�͂�c�uD�Y#5>�X<�i	e
��i�d�8�!��h��+^O�q���GR�)$��P�;��)��02���{��x�u�S�G�����Ê��k�kY�#���dfbF�U�ir x���\��3��q4�����Ud%�6,�X�s��h�:����p�#llY��	��h�F��ުJ��H��s���ג�
�{)&y�h�0��L �^p��cĮ_��L���m�B��"����feB4Đ�X��Ǫ/�9æ����a� >j)��_o��`������R&u�Լ܎<G�1.���*��F�F
�YB2�؃����89��\׸hS�c�ph�U�Yu��9�B��h�#�R�c��MfY�R�����>Qv4�F��	c� �c�׿X�'D[[��/+@����C=��ϰ#�P[z��z}�SC��&T��C�jI�s1G_��$����L�z�(��5��Tqٰ")��(��J�:����m q���"O�dwhfmm�����-�|ߍ��TN���p�rV�Б9D�ڨaj�n���F��
���Ff�
�  �H\o�X7'A<�me�Ju��}H\3V�D\��$n�e�&lI���`�G�Uy^V�Wܮ�T�� �c��W�ER�e�j�Q�ro -�A�'*yi��T'�����?���k���SF~py�rЇ��N��!Txח4`��Z����nض�Ђ>��i��v.��T�!.�X�i��Hl^r��	�s���'�Y�R@�UƔ.Yr�a:�ж3�>i�K3\��1��~]�]_�����V4_��S
�W������.S�,��.]�
�ҤH����r�����s�*��=sw)��1PI�:�۷������2UY�eק���p�{z���K���r%�H���M~3��R�4P�}�m�c0�d�D��Vˈ�Wp����ml�*�ܚq�w�,~r��#ilUǮ������p�,)�4S��c��ߚ��5#�K�3�����"pX����1�����-�ܿ`_x4Ϭ���6���g����s[G��B�ĴP�xR���EǞZR�ʕ� �C���j� �v�>�ZecD��g�
΍�Z\���;9P�{��)�tCU+���_t�́��1����38��Z�X��@�욬5zoF |�
�r�{- ���a�Y�<��k��_1�ki�!"1"���&^B�uXȍ"E��0`���2��5���ʞ���=��k���m������F�iX�T#���HYE��U,2��`U���E���ĳ�9�`��h��U.n| {�C�@�d\J{!?:��`F���N��B��������D� Ί_��=��۾�Cd}ې��V?f�q�d��N����I?EM]v��*D}�h�RRЩ;x$�`��Fg:H����w�V������*_�9'�yY�r�|��n���U���ޡ�3f�)� ��f�G�U�(���LI��0�+ޓA���X{+���W8W�ji��a�,ڂ�-�-�p���"��`���3��s�"l9��ܪ���m�b�kX��	���j��8I�79Tq��*���s�Hy�0r5 _��J���7z�>��R*P��
�+E�?o�q3���x߅��`py��E�k���2�T�j5(�,rI����Y8�l�*���@釠���6��+��3�UT9��WhjL�U����Rq����[�^a�%�݆9��09D�f^�����#����FނxY#���o���98������d��$�W�bĬ����W'/,�rs���l�6��W ��!V�z?�T�J�1�9.w��H�I��d8�8����&���JTͥ�ވ���+�Ɩ��G���eK��*uZ:�A�@�-o�(F�YG�#=����7�H:4?��MtBb��<���|�9�*7v�S�
�$w�u�xCp�����W�L�&�H8�l.�1��O�>��uj�!�t��銏������.����}?�dJ�9k�>�S��H��F�K�8���Q�2����dOp!�c�-�� L\�ĺ�:S��_w����n7*@��C_ЊL�Y��� 	>܁<��뀽�X2��N�����e��m�oR*�KM��V(�ul�W�tQNO��3���K��;5FZ�Iw�D��a�wr��R���3Y���َX��I�� �c��yfv������>v�P�o7�Pz{D��g�/i��<���Ğp�����P8|h�<b�}4�y\+�q�n&*�W�1Jqt	@�V~�*,�����tu�֑��Ծ wK�gA�GM���Xj=S�:5��U>�긴�c%�+?��'�<��`Ȉ��~�Ci�y6�m�mȒ��fF 9���P��H�t����҄�p��(��ud썊4�'���G#0�IV�	M	�_c�#�EFJ� ۫i�D��!;lx�.ϗ�_�fD����e@�=����p��Ho�=h���&R��1!� �Y����E�<�vZ����Z�ºQ(Cv[�Dy���������H�ϻX�-.��#rs���2v<���	��v��9���	��m�MB�N���H<Ҍ�1P�����~��(��|�V=[#���z��L�����ݮ��8?*�"9���1l���?�"w���c�W-%���	{V"�Q�C���o��V��ȑ`��9�CC�b΢M��4�4M�ɣ�#��
�GP�����t��:��{�dw@F Ts��`gM{�6�&5�&	���E�8�Y.�ڦ�=�ɞ�E��
\�#C?~'<�B��
ya��i��Ik���8��<�|�$��1���f�F#�a���7�1����Q�x�$�fF`��%F�f��K���;t#�P�>����|؎ɨc�T���6F3g��6���'������� d-���Z�5��y9hw��Z�i7uh��<(�o}F} �wfS�)���;���'���д�j�����F��=�vK�c~��U�\kS��W��o<Ŧ������$�+k�GGo]�^�Q{EO��fx�ЗTm%��Pj���O��A����%�3�^#wF�ߞg�1���KL,B�j
1�E2z눊�SS�%dt�.EW��h0�Λ���@�LuZ�7�e�E<Mj�Yy��|�<��\nu��M�\m9k�`��J/��t�+9�����/2f�y~�@vߢE�"Xژ'i�54�=ii4;O�-[�w���zױ�����③r�d���\��ꮈ3ќ�˞/��J�8����G\���CF�;F���11��UۼH�];�%I��l���y���J�I��)��3�E[h8��M��&BT�K�&�Uz�"��2̓y�1�� L� �.��*��LƆYܝ���c3B��.}����e\�2�:�jgQ��?9A���'k��:��B�Qz�H��=�T������H��.#:�����Ғ�����j��s����#���*$�/r��
�d����ܲx�<Y�kv1�t8\4�gC�3�ձ�z�f}��a�-� ���JL~m���GҁBk��u�Dd�~��}���Т�c�0w���cqZ,`8����ܓ$:�+�&�95)dp�H�I,GF3R�ka/&��"���6ˌ<�T<��"���Y���b�e�c|�� $��X��O�M���&����L��>��xra{��#�V=�B6���i���ǻ��DI�_���K��d����wߘXB@�R?�Ȯ>ө8&� ���
g�[�;#�?N{G�����<���A4��j-:&1.���M?��@�r���2�����\P9+|���>�q���]Ա����
���������[������\�=U(���5\lB���!��C��&^�.���<I�6��^�vY�����4}.ԝ
Ȏ�����
�~.�L�q0��C�+Ա>��Ɏ�-�S��?�|V��,��tT?��}�}�0w��=0��
y�0�ߝ$�
������컆��������16A���(�l��e���Z��/�S2_j���l,���	(r����k @d��h[��W�<����'�R�D;Mt$^��#��g��