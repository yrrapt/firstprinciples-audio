XlxV65EB     d38     400sgӮ�,�W�u��*���>��ߌH��څC;�W!w[�&���Ь\p��yYnp���2��G�LQ���a?J�*����,�M��4� >���?L;���fx���y��n���k�o�Eqr�O�a�Fq��
���2�hZ�3	Ժ�'���y�3%�o�\�NG��d8��|ݖ��s
5�y��)���� U+^p�K�*(Q�4���|�	��G#��e	 �T!J�k`?��1[��o>|Y��&�;qY���q��d!Hie&���ط��1a��8�����I�':R��`����wao��A��ژ媏���F�9?�z��.*����.�����ن��NlMhޝ�mq�(s��V����"��,͌,�8[�s���� ���P��G�A��~n���"�×���*�=���7^`�}�Z�%r�/)�%��ޱ#&�d��_����M�V�g�d�����NJ5G~V�[�1�֦2���'G$i"e0Y;���.�ϮrCtm㽎=U*.�~���7���[�JM;'rԆ�y6po�M�i��"��E�a�V��n�D�iڕ͗�F�̡�_?cҦAm�F��&B����ȭ���n7�����A���'m�կ��
�]�yv
dh6GX�;��ڦ���p@�#�<���^eES�j�YT�NІ�,U��?���{j$N{��m"Bs����q��ؾI��̉4��#kl�f��Š�\?�.���ie;����� �"P�4Ag�n��)�/�f*�mwR`��0��mI�\9�\Ct��s&+�X1"tcDX��W(#4����|�``��Ơ��s��H��J�G��K^�����7��Ba>�����2Axk�t���/���
$���NQ���'��L�!�9�(���U��%s��ó�5�.1EhVG�����b���Z,/��܏��"�v��xm�gL�v��ƟЕ��opw��FĪ�H��	A�h_lR�t�$�y .��c�:9������4��9�